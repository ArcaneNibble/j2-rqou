-- Copyright (c) 2015, Smart Energy Instruments Inc.
-- All rights reserved.  For details, see COPYING in the top level directory.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package attr_pack is

  -- There is a global namespace for connecting signals and ports within a
  -- design. The soc_gen tool will connect ports with matching names. If a port
  -- is insided a global_ports group, its port name becomes it's global signal
  -- name. An sei_port_global_name attribute explicitly sets a ports global
  -- name to something different than the port name.
  -- A port can have a local name, in which case it's global name will
  -- generated by prefixing the global name with the device's name. A
  -- device named "dev0" with a local port "rx" will have the rx port connected
  -- to the global signal "dev0_rx". Like global ports, the name of a local
  -- port can be overridden by an attribute, sei_port_local_name.

-- synopsys translate_off
  -- groups entity ports that are local ports. They will be connected in the
  -- global namespace, but their name is first prefixed by the device name. Use
  -- sei_port_local_name instead to override the port name.
  group local_ports is (signal <>);
  -- groups entity ports that are global ports. They will be connected in the
  -- global namespace using the port's name. Use sei_port_global_name instead
  -- to override the port name.
  group global_ports is (signal <>);
  -- groups ports that connecting to the ring bus
  group bus_ports is (signal <>);
-- synopsys translate_on

  -- sets the global name of a port
  attribute sei_port_global_name : string;
  -- sets the local name of a port
  attribute sei_port_local_name : string;

  -- identify entity ports that are clocks
  attribute sei_port_clock : boolean;

  -- identify entity port that is an irq line
  attribute sei_port_irq : boolean;

  -- name of the target technology that an architecture is suited for
  -- eg. "spartan6", "kintex7", "tsmc"
  attribute sei_target : string;
end package;
