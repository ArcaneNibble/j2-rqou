library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.sgs1010d_pack.all;

entity digitial_top_tb is
end digital_top_tb;

architecture tb of digital_top_tb is
begin

end tb;
